type rom_array is array (natural range <>) of std_logic_vector ( 63 downto 0 ) ;
constant  rom : rom_array := ( 
--  Master code
 x"0c00_0000_0018_ffff", -- 0
 x"8002_201f_a402_1400", -- 4
 x"2001_a003_400f_6000", -- 8
 x"8812_c820_81fa_8812", -- c
 x"c820_1000_0000_0004", -- 10
 x"2000_a003_1400_ffff", -- 14
 x"1000_0000_0008_1c00", -- 18
 x"ffff_ffff_ffff_ffff", -- 1c
--  Slave code
 x"1000_0000_0040_1c00", -- 0
 x"c814_8a02_2001_c836", -- 4
 x"a000_0403_8810_a000", -- 8
 x"1400_ffff_ffff_ffff", -- c
 x"2000_2000_2008_c82d", -- 10
 x"2000_a007_a007_8810", -- 14
 x"a000_8810_b008_2fff", -- 18
 x"c825_d009_2014_c82b", -- 1c
 x"2fff_c825_b008_c814", -- 20
 x"d009_b008_c814_c820", -- 24
 x"2001_2ffe_c82d_c83c", -- 28
 x"a000_0403_a822_ffff", -- 2c
 x"8806_a823_8007_a833", -- 30
 x"a000_07e2_8006_8006", -- 34
 x"a201_1400_ffff_ffff", -- 38
 x"1000_0000_0010_1c00", -- 3c
 x"1000_0000_0005_1400", -- 40
 x"ffff_ffff_ffff_ffff"  -- 44
);
